// Copyright 2022 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// FPU Subsystem Instruction Package
// Contributor: Fabio Cappellini <fcappellini@ethz.ch>


  package fpu_ss_instr_pkg;

  localparam logic [15:0] C_FLWSP            = 16'b011???????????10;
  localparam logic [15:0] C_FSWSP            = 16'b111???????????10;
  localparam logic [15:0] C_FLW              = 16'b011???????????00;
  localparam logic [15:0] C_FSW              = 16'b111???????????00;


  localparam logic [31:0] CSRRW_FSCSR        = 32'b000000000011?????001?????1110011;
  localparam logic [31:0] CSRRS_FRCSR        = 32'b000000000011?????010?????1110011;
  localparam logic [31:0] CSRRW_FSRM         = 32'b000000000010?????001?????1110011;
  localparam logic [31:0] CSRRS_FRRM         = 32'b000000000010?????010?????1110011;
  localparam logic [31:0] CSRRWI_FSRMI       = 32'b000000000010?????101?????1110011;
  localparam logic [31:0] CSRRW_FSFLAGS      = 32'b000000000001?????001?????1110011;
  localparam logic [31:0] CSRRS_FRFLAGS      = 32'b000000000001?????010?????1110011;
  localparam logic [31:0] CSRRWI_FSFLAGSI    = 32'b000000000001?????101?????1110011;

  localparam logic [31:0] CSRRW_FSMODE       = 32'b100000000000?????001?????1110011;
  localparam logic [31:0] CSRRS_FRMODE       = 32'b100000000000?????010?????1110011;
  localparam logic [31:0] CSRRWI_FSMODEI     = 32'b100000000000?????101?????1110011;

  localparam logic [31:0] CSRRW_FSSRM        = 32'b100000000001?????001?????1110011;
  localparam logic [31:0] CSRRS_FRSRM        = 32'b100000000001?????010?????1110011;
  localparam logic [31:0] CSRRWI_FSSRMI      = 32'b100000000001?????101?????1110011;


  localparam logic [31:0] BEQ                = 32'b?????????????????000?????1100011;
  localparam logic [31:0] BNE                = 32'b?????????????????001?????1100011;
  localparam logic [31:0] BLT                = 32'b?????????????????100?????1100011;
  localparam logic [31:0] BGE                = 32'b?????????????????101?????1100011;
  localparam logic [31:0] BLTU               = 32'b?????????????????110?????1100011;
  localparam logic [31:0] BGEU               = 32'b?????????????????111?????1100011;
  localparam logic [31:0] JALR               = 32'b?????????????????000?????1100111;
  localparam logic [31:0] JAL                = 32'b?????????????????????????1101111;
  localparam logic [31:0] LUI                = 32'b?????????????????????????0110111;
  localparam logic [31:0] AUIPC              = 32'b?????????????????????????0010111;
  localparam logic [31:0] ADDI               = 32'b?????????????????000?????0010011;
  localparam logic [31:0] SLLI               = 32'b000000???????????001?????0010011;
  localparam logic [31:0] SLTI               = 32'b?????????????????010?????0010011;
  localparam logic [31:0] SLTIU              = 32'b?????????????????011?????0010011;
  localparam logic [31:0] XORI               = 32'b?????????????????100?????0010011;
  localparam logic [31:0] SRLI               = 32'b000000???????????101?????0010011;
  localparam logic [31:0] SRAI               = 32'b010000???????????101?????0010011;
  localparam logic [31:0] ORI                = 32'b?????????????????110?????0010011;
  localparam logic [31:0] ANDI               = 32'b?????????????????111?????0010011;
  localparam logic [31:0] ADD                = 32'b0000000??????????000?????0110011;
  localparam logic [31:0] SUB                = 32'b0100000??????????000?????0110011;
  localparam logic [31:0] SLL                = 32'b0000000??????????001?????0110011;
  localparam logic [31:0] SLT                = 32'b0000000??????????010?????0110011;
  localparam logic [31:0] SLTU               = 32'b0000000??????????011?????0110011;
  localparam logic [31:0] XOR                = 32'b0000000??????????100?????0110011;
  localparam logic [31:0] SRL                = 32'b0000000??????????101?????0110011;
  localparam logic [31:0] SRA                = 32'b0100000??????????101?????0110011;
  localparam logic [31:0] OR                 = 32'b0000000??????????110?????0110011;
  localparam logic [31:0] AND                = 32'b0000000??????????111?????0110011;
  localparam logic [31:0] ADDIW              = 32'b?????????????????000?????0011011;
  localparam logic [31:0] SLLIW              = 32'b0000000??????????001?????0011011;
  localparam logic [31:0] SRLIW              = 32'b0000000??????????101?????0011011;
  localparam logic [31:0] SRAIW              = 32'b0100000??????????101?????0011011;
  localparam logic [31:0] ADDW               = 32'b0000000??????????000?????0111011;
  localparam logic [31:0] SUBW               = 32'b0100000??????????000?????0111011;
  localparam logic [31:0] SLLW               = 32'b0000000??????????001?????0111011;
  localparam logic [31:0] SRLW               = 32'b0000000??????????101?????0111011;
  localparam logic [31:0] SRAW               = 32'b0100000??????????101?????0111011;
  localparam logic [31:0] LB                 = 32'b?????????????????000?????0000011;
  localparam logic [31:0] LH                 = 32'b?????????????????001?????0000011;
  localparam logic [31:0] LW                 = 32'b?????????????????010?????0000011;
  localparam logic [31:0] LD                 = 32'b?????????????????011?????0000011;
  localparam logic [31:0] LBU                = 32'b?????????????????100?????0000011;
  localparam logic [31:0] LHU                = 32'b?????????????????101?????0000011;
  localparam logic [31:0] LWU                = 32'b?????????????????110?????0000011;
  localparam logic [31:0] SB                 = 32'b?????????????????000?????0100011;
  localparam logic [31:0] SH                 = 32'b?????????????????001?????0100011;
  localparam logic [31:0] SW                 = 32'b?????????????????010?????0100011;
  localparam logic [31:0] SD                 = 32'b?????????????????011?????0100011;
  localparam logic [31:0] FENCE              = 32'b?????????????????000?????0001111;
  localparam logic [31:0] FENCE_I            = 32'b?????????????????001?????0001111;
  localparam logic [31:0] MUL                = 32'b0000001??????????000?????0110011;
  localparam logic [31:0] MULH               = 32'b0000001??????????001?????0110011;
  localparam logic [31:0] MULHSU             = 32'b0000001??????????010?????0110011;
  localparam logic [31:0] MULHU              = 32'b0000001??????????011?????0110011;
  localparam logic [31:0] DIV                = 32'b0000001??????????100?????0110011;
  localparam logic [31:0] DIVU               = 32'b0000001??????????101?????0110011;
  localparam logic [31:0] REM                = 32'b0000001??????????110?????0110011;
  localparam logic [31:0] REMU               = 32'b0000001??????????111?????0110011;
  localparam logic [31:0] MULW               = 32'b0000001??????????000?????0111011;
  localparam logic [31:0] DIVW               = 32'b0000001??????????100?????0111011;
  localparam logic [31:0] DIVUW              = 32'b0000001??????????101?????0111011;
  localparam logic [31:0] REMW               = 32'b0000001??????????110?????0111011;
  localparam logic [31:0] REMUW              = 32'b0000001??????????111?????0111011;
  localparam logic [31:0] ANDN               = 32'b0100000??????????111?????0110011;
  localparam logic [31:0] ORN                = 32'b0100000??????????110?????0110011;
  localparam logic [31:0] XNOR               = 32'b0100000??????????100?????0110011;
  localparam logic [31:0] SLO                = 32'b0010000??????????001?????0110011;
  localparam logic [31:0] SRO                = 32'b0010000??????????101?????0110011;
  localparam logic [31:0] ROL                = 32'b0110000??????????001?????0110011;
  localparam logic [31:0] ROR                = 32'b0110000??????????101?????0110011;
  localparam logic [31:0] SBCLR              = 32'b0100100??????????001?????0110011;
  localparam logic [31:0] SBSET              = 32'b0010100??????????001?????0110011;
  localparam logic [31:0] SBINV              = 32'b0110100??????????001?????0110011;
  localparam logic [31:0] SBEXT              = 32'b0100100??????????101?????0110011;
  localparam logic [31:0] GORC               = 32'b0010100??????????101?????0110011;
  localparam logic [31:0] GREV               = 32'b0110100??????????101?????0110011;
  localparam logic [31:0] SLOI               = 32'b001000???????????001?????0010011;
  localparam logic [31:0] SROI               = 32'b001000???????????101?????0010011;
  localparam logic [31:0] RORI               = 32'b011000???????????101?????0010011;
  localparam logic [31:0] SBCLRI             = 32'b010010???????????001?????0010011;
  localparam logic [31:0] SBSETI             = 32'b001010???????????001?????0010011;
  localparam logic [31:0] SBINVI             = 32'b011010???????????001?????0010011;
  localparam logic [31:0] SBEXTI             = 32'b010010???????????101?????0010011;
  localparam logic [31:0] GORCI              = 32'b001010???????????101?????0010011;
  localparam logic [31:0] GREVI              = 32'b011010???????????101?????0010011;
  localparam logic [31:0] CMIX               = 32'b?????11??????????001?????0110011;
  localparam logic [31:0] CMOV               = 32'b?????11??????????101?????0110011;
  localparam logic [31:0] FSL                = 32'b?????10??????????001?????0110011;
  localparam logic [31:0] FSR                = 32'b?????10??????????101?????0110011;
  localparam logic [31:0] FSRI               = 32'b?????1???????????101?????0010011;
  localparam logic [31:0] CLZ                = 32'b011000000000?????001?????0010011;
  localparam logic [31:0] CTZ                = 32'b011000000001?????001?????0010011;
  localparam logic [31:0] PCNT               = 32'b011000000010?????001?????0010011;
  localparam logic [31:0] SEXT_B             = 32'b011000000100?????001?????0010011;
  localparam logic [31:0] SEXT_H             = 32'b011000000101?????001?????0010011;
  localparam logic [31:0] CRC32_B            = 32'b011000010000?????001?????0010011;
  localparam logic [31:0] CRC32_H            = 32'b011000010001?????001?????0010011;
  localparam logic [31:0] CRC32_W            = 32'b011000010010?????001?????0010011;
  localparam logic [31:0] CRC32C_B           = 32'b011000011000?????001?????0010011;
  localparam logic [31:0] CRC32C_H           = 32'b011000011001?????001?????0010011;
  localparam logic [31:0] CRC32C_W           = 32'b011000011010?????001?????0010011;
  localparam logic [31:0] SH1ADD             = 32'b0010000??????????010?????0110011;
  localparam logic [31:0] SH2ADD             = 32'b0010000??????????100?????0110011;
  localparam logic [31:0] SH3ADD             = 32'b0010000??????????110?????0110011;
  localparam logic [31:0] CLMUL              = 32'b0000101??????????001?????0110011;
  localparam logic [31:0] CLMULR             = 32'b0000101??????????010?????0110011;
  localparam logic [31:0] CLMULH             = 32'b0000101??????????011?????0110011;
  localparam logic [31:0] MIN                = 32'b0000101??????????100?????0110011;
  localparam logic [31:0] MAX                = 32'b0000101??????????101?????0110011;
  localparam logic [31:0] MINU               = 32'b0000101??????????110?????0110011;
  localparam logic [31:0] MAXU               = 32'b0000101??????????111?????0110011;
  localparam logic [31:0] SHFL               = 32'b0000100??????????001?????0110011;
  localparam logic [31:0] UNSHFL             = 32'b0000100??????????101?????0110011;
  localparam logic [31:0] BEXT               = 32'b0000100??????????110?????0110011;
  localparam logic [31:0] BDEP               = 32'b0100100??????????110?????0110011;
  localparam logic [31:0] PACK               = 32'b0000100??????????100?????0110011;
  localparam logic [31:0] PACKU              = 32'b0100100??????????100?????0110011;
  localparam logic [31:0] PACKH              = 32'b0000100??????????111?????0110011;
  localparam logic [31:0] BFP                = 32'b0100100??????????111?????0110011;
  localparam logic [31:0] SHFLI              = 32'b0000100??????????001?????0010011;
  localparam logic [31:0] UNSHFLI            = 32'b0000100??????????101?????0010011;
  localparam logic [31:0] AMOADD_W           = 32'b00000????????????010?????0101111;
  localparam logic [31:0] AMOXOR_W           = 32'b00100????????????010?????0101111;
  localparam logic [31:0] AMOOR_W            = 32'b01000????????????010?????0101111;
  localparam logic [31:0] AMOAND_W           = 32'b01100????????????010?????0101111;
  localparam logic [31:0] AMOMIN_W           = 32'b10000????????????010?????0101111;
  localparam logic [31:0] AMOMAX_W           = 32'b10100????????????010?????0101111;
  localparam logic [31:0] AMOMINU_W          = 32'b11000????????????010?????0101111;
  localparam logic [31:0] AMOMAXU_W          = 32'b11100????????????010?????0101111;
  localparam logic [31:0] AMOSWAP_W          = 32'b00001????????????010?????0101111;
  localparam logic [31:0] LR_W               = 32'b00010??00000?????010?????0101111;
  localparam logic [31:0] SC_W               = 32'b00011????????????010?????0101111;
  localparam logic [31:0] AMOADD_D           = 32'b00000????????????011?????0101111;
  localparam logic [31:0] AMOXOR_D           = 32'b00100????????????011?????0101111;
  localparam logic [31:0] AMOOR_D            = 32'b01000????????????011?????0101111;
  localparam logic [31:0] AMOAND_D           = 32'b01100????????????011?????0101111;
  localparam logic [31:0] AMOMIN_D           = 32'b10000????????????011?????0101111;
  localparam logic [31:0] AMOMAX_D           = 32'b10100????????????011?????0101111;
  localparam logic [31:0] AMOMINU_D          = 32'b11000????????????011?????0101111;
  localparam logic [31:0] AMOMAXU_D          = 32'b11100????????????011?????0101111;
  localparam logic [31:0] AMOSWAP_D          = 32'b00001????????????011?????0101111;
  localparam logic [31:0] LR_D               = 32'b00010??00000?????011?????0101111;
  localparam logic [31:0] SC_D               = 32'b00011????????????011?????0101111;
  localparam logic [31:0] ECALL              = 32'b00000000000000000000000001110011;
  localparam logic [31:0] EBREAK             = 32'b00000000000100000000000001110011;
  localparam logic [31:0] URET               = 32'b00000000001000000000000001110011;
  localparam logic [31:0] SRET               = 32'b00010000001000000000000001110011;
  localparam logic [31:0] MRET               = 32'b00110000001000000000000001110011;
  localparam logic [31:0] DRET               = 32'b01111011001000000000000001110011;
  localparam logic [31:0] SFENCE_VMA         = 32'b0001001??????????000000001110011;
  localparam logic [31:0] WFI                = 32'b00010000010100000000000001110011;
  localparam logic [31:0] CSRRW              = 32'b?????????????????001?????1110011;
  localparam logic [31:0] CSRRS              = 32'b?????????????????010?????1110011;
  localparam logic [31:0] CSRRC              = 32'b?????????????????011?????1110011;
  localparam logic [31:0] CSRRWI             = 32'b?????????????????101?????1110011;
  localparam logic [31:0] CSRRSI             = 32'b?????????????????110?????1110011;
  localparam logic [31:0] CSRRCI             = 32'b?????????????????111?????1110011;
  localparam logic [31:0] HFENCE_BVMA        = 32'b0010001??????????000000001110011;
  localparam logic [31:0] HFENCE_GVMA        = 32'b1010001??????????000000001110011;
  localparam logic [31:0] FADD_S             = 32'b0000000??????????????????1010011;
  localparam logic [31:0] FSUB_S             = 32'b0000100??????????????????1010011;
  localparam logic [31:0] FMUL_S             = 32'b0001000??????????????????1010011;
  localparam logic [31:0] FDIV_S             = 32'b0001100??????????????????1010011;
  localparam logic [31:0] FSGNJ_S            = 32'b0010000??????????000?????1010011;
  localparam logic [31:0] FSGNJN_S           = 32'b0010000??????????001?????1010011;
  localparam logic [31:0] FSGNJX_S           = 32'b0010000??????????010?????1010011;
  localparam logic [31:0] FMIN_S             = 32'b0010100??????????000?????1010011;
  localparam logic [31:0] FMAX_S             = 32'b0010100??????????001?????1010011;
  localparam logic [31:0] FSQRT_S            = 32'b010110000000?????????????1010011;
  localparam logic [31:0] FADD_D             = 32'b0000001??????????????????1010011;
  localparam logic [31:0] FSUB_D             = 32'b0000101??????????????????1010011;
  localparam logic [31:0] FMUL_D             = 32'b0001001??????????????????1010011;
  localparam logic [31:0] FDIV_D             = 32'b0001101??????????????????1010011;
  localparam logic [31:0] FSGNJ_D            = 32'b0010001??????????000?????1010011;
  localparam logic [31:0] FSGNJN_D           = 32'b0010001??????????001?????1010011;
  localparam logic [31:0] FSGNJX_D           = 32'b0010001??????????010?????1010011;
  localparam logic [31:0] FMIN_D             = 32'b0010101??????????000?????1010011;
  localparam logic [31:0] FMAX_D             = 32'b0010101??????????001?????1010011;
  localparam logic [31:0] FCVT_S_D           = 32'b010000000001?????????????1010011;
  localparam logic [31:0] FCVT_D_S           = 32'b010000100000?????????????1010011;
  localparam logic [31:0] FSQRT_D            = 32'b010110100000?????????????1010011;
  localparam logic [31:0] FADD_Q             = 32'b0000011??????????????????1010011;
  localparam logic [31:0] FSUB_Q             = 32'b0000111??????????????????1010011;
  localparam logic [31:0] FMUL_Q             = 32'b0001011??????????????????1010011;
  localparam logic [31:0] FDIV_Q             = 32'b0001111??????????????????1010011;
  localparam logic [31:0] FSGNJ_Q            = 32'b0010011??????????000?????1010011;
  localparam logic [31:0] FSGNJN_Q           = 32'b0010011??????????001?????1010011;
  localparam logic [31:0] FSGNJX_Q           = 32'b0010011??????????010?????1010011;
  localparam logic [31:0] FMIN_Q             = 32'b0010111??????????000?????1010011;
  localparam logic [31:0] FMAX_Q             = 32'b0010111??????????001?????1010011;
  localparam logic [31:0] FCVT_S_Q           = 32'b010000000011?????????????1010011;
  localparam logic [31:0] FCVT_Q_S           = 32'b010001100000?????????????1010011;
  localparam logic [31:0] FCVT_D_Q           = 32'b010000100011?????????????1010011;
  localparam logic [31:0] FCVT_Q_D           = 32'b010001100001?????????????1010011;
  localparam logic [31:0] FSQRT_Q            = 32'b010111100000?????????????1010011;
  localparam logic [31:0] FLE_S              = 32'b1010000??????????000?????1010011;
  localparam logic [31:0] FLT_S              = 32'b1010000??????????001?????1010011;
  localparam logic [31:0] FEQ_S              = 32'b1010000??????????010?????1010011;
  localparam logic [31:0] FLE_D              = 32'b1010001??????????000?????1010011;
  localparam logic [31:0] FLT_D              = 32'b1010001??????????001?????1010011;
  localparam logic [31:0] FEQ_D              = 32'b1010001??????????010?????1010011;
  localparam logic [31:0] FLE_Q              = 32'b1010011??????????000?????1010011;
  localparam logic [31:0] FLT_Q              = 32'b1010011??????????001?????1010011;
  localparam logic [31:0] FEQ_Q              = 32'b1010011??????????010?????1010011;
  localparam logic [31:0] FCVT_W_S           = 32'b110000000000?????????????1010011;
  localparam logic [31:0] FCVT_WU_S          = 32'b110000000001?????????????1010011;
  localparam logic [31:0] FCVT_L_S           = 32'b110000000010?????????????1010011;
  localparam logic [31:0] FCVT_LU_S          = 32'b110000000011?????????????1010011;
  localparam logic [31:0] FMV_X_W            = 32'b111000000000?????000?????1010011;
  localparam logic [31:0] FCLASS_S           = 32'b111000000000?????001?????1010011;
  localparam logic [31:0] FCVT_W_D           = 32'b110000100000?????????????1010011;
  localparam logic [31:0] FCVT_WU_D          = 32'b110000100001?????????????1010011;
  localparam logic [31:0] FCVT_L_D           = 32'b110000100010?????????????1010011;
  localparam logic [31:0] FCVT_LU_D          = 32'b110000100011?????????????1010011;
  localparam logic [31:0] FMV_X_D            = 32'b111000100000?????000?????1010011;
  localparam logic [31:0] FCLASS_D           = 32'b111000100000?????001?????1010011;
  localparam logic [31:0] FCVT_W_Q           = 32'b110001100000?????????????1010011;
  localparam logic [31:0] FCVT_WU_Q          = 32'b110001100001?????????????1010011;
  localparam logic [31:0] FCVT_L_Q           = 32'b110001100010?????????????1010011;
  localparam logic [31:0] FCVT_LU_Q          = 32'b110001100011?????????????1010011;
  localparam logic [31:0] FMV_X_Q            = 32'b111001100000?????000?????1010011;
  localparam logic [31:0] FCLASS_Q           = 32'b111001100000?????001?????1010011;
  localparam logic [31:0] FCVT_S_W           = 32'b110100000000?????????????1010011;
  localparam logic [31:0] FCVT_S_WU          = 32'b110100000001?????????????1010011;
  localparam logic [31:0] FCVT_S_L           = 32'b110100000010?????????????1010011;
  localparam logic [31:0] FCVT_S_LU          = 32'b110100000011?????????????1010011;
  localparam logic [31:0] FMV_W_X            = 32'b111100000000?????000?????1010011;
  localparam logic [31:0] FCVT_D_W           = 32'b110100100000?????????????1010011;
  localparam logic [31:0] FCVT_D_WU          = 32'b110100100001?????????????1010011;
  localparam logic [31:0] FCVT_D_L           = 32'b110100100010?????????????1010011;
  localparam logic [31:0] FCVT_D_LU          = 32'b110100100011?????????????1010011;
  localparam logic [31:0] FMV_D_X            = 32'b111100100000?????000?????1010011;
  localparam logic [31:0] FCVT_Q_W           = 32'b110101100000?????????????1010011;
  localparam logic [31:0] FCVT_Q_WU          = 32'b110101100001?????????????1010011;
  localparam logic [31:0] FCVT_Q_L           = 32'b110101100010?????????????1010011;
  localparam logic [31:0] FCVT_Q_LU          = 32'b110101100011?????????????1010011;
  localparam logic [31:0] FMV_Q_X            = 32'b111101100000?????000?????1010011;
  localparam logic [31:0] FLW                = 32'b?????????????????010?????0000111;
  localparam logic [31:0] FLD                = 32'b?????????????????011?????0000111;
  localparam logic [31:0] FLQ                = 32'b?????????????????100?????0000111;
  localparam logic [31:0] FSW                = 32'b?????????????????010?????0100111;
  localparam logic [31:0] FSD                = 32'b?????????????????011?????0100111;
  localparam logic [31:0] FSQ                = 32'b?????????????????100?????0100111;
  localparam logic [31:0] FMADD_S            = 32'b?????00??????????????????1000011;
  localparam logic [31:0] FMSUB_S            = 32'b?????00??????????????????1000111;
  localparam logic [31:0] FNMSUB_S           = 32'b?????00??????????????????1001011;
  localparam logic [31:0] FNMADD_S           = 32'b?????00??????????????????1001111;
  localparam logic [31:0] FMADD_D            = 32'b?????01??????????????????1000011;
  localparam logic [31:0] FMSUB_D            = 32'b?????01??????????????????1000111;
  localparam logic [31:0] FNMSUB_D           = 32'b?????01??????????????????1001011;
  localparam logic [31:0] FNMADD_D           = 32'b?????01??????????????????1001111;
  localparam logic [31:0] FMADD_Q            = 32'b?????11??????????????????1000011;
  localparam logic [31:0] FMSUB_Q            = 32'b?????11??????????????????1000111;
  localparam logic [31:0] FNMSUB_Q           = 32'b?????11??????????????????1001011;
  localparam logic [31:0] FNMADD_Q           = 32'b?????11??????????????????1001111;
  localparam logic [31:0] DMSRC              = 32'b0000000??????????000000000101011;
  localparam logic [31:0] DMDST              = 32'b0000001??????????000000000101011;
  localparam logic [31:0] DMCPYI             = 32'b0000010??????????000?????0101011;
  localparam logic [31:0] DMCPY              = 32'b0000011??????????000?????0101011;
  localparam logic [31:0] DMSTATI            = 32'b0000100?????00000000?????0101011;
  localparam logic [31:0] DMSTAT             = 32'b0000101?????00000000?????0101011;
  localparam logic [31:0] DMSTR              = 32'b0000110??????????000000000101011;
  localparam logic [31:0] DMREP              = 32'b000011100000?????000000000101011;
  localparam logic [31:0] FREP_O             = 32'b????????????????????????10001011;
  localparam logic [31:0] FREP_I             = 32'b????????????????????????00001011;
  localparam logic [31:0] IREP               = 32'b?????????????????????????0111111;
  localparam logic [31:0] SCFGRI             = 32'b????????????00000001?????0101011;
  localparam logic [31:0] SCFGWI             = 32'b?????????????????010000000101011;
  localparam logic [31:0] SCFGR              = 32'b0000000?????00001001?????0101011;
  localparam logic [31:0] SCFGW              = 32'b0000000??????????010000010101011;
  localparam logic [31:0] FLH                = 32'b?????????????????001?????0000111;
  localparam logic [31:0] FSH                = 32'b?????????????????001?????0100111;
  localparam logic [31:0] FMADD_H            = 32'b?????10??????????????????1000011;
  localparam logic [31:0] FMSUB_H            = 32'b?????10??????????????????1000111;
  localparam logic [31:0] FNMSUB_H           = 32'b?????10??????????????????1001011;
  localparam logic [31:0] FNMADD_H           = 32'b?????10??????????????????1001111;
  localparam logic [31:0] FADD_H             = 32'b0000010??????????????????1010011;
  localparam logic [31:0] FSUB_H             = 32'b0000110??????????????????1010011;
  localparam logic [31:0] FMUL_H             = 32'b0001010??????????????????1010011;
  localparam logic [31:0] FDIV_H             = 32'b0001110??????????????????1010011;
  localparam logic [31:0] FSQRT_H            = 32'b010111000000?????????????1010011;
  localparam logic [31:0] FSGNJ_H            = 32'b0010010??????????000?????1010011;
  localparam logic [31:0] FSGNJN_H           = 32'b0010010??????????001?????1010011;
  localparam logic [31:0] FSGNJX_H           = 32'b0010010??????????010?????1010011;
  localparam logic [31:0] FMIN_H             = 32'b0010110??????????000?????1010011;
  localparam logic [31:0] FMAX_H             = 32'b0010110??????????001?????1010011;
  localparam logic [31:0] FEQ_H              = 32'b1010010??????????010?????1010011;
  localparam logic [31:0] FLT_H              = 32'b1010010??????????001?????1010011;
  localparam logic [31:0] FLE_H              = 32'b1010010??????????000?????1010011;
  localparam logic [31:0] FCVT_W_H           = 32'b110001000000?????????????1010011;
  localparam logic [31:0] FCVT_WU_H          = 32'b110001000001?????????????1010011;
  localparam logic [31:0] FCVT_H_W           = 32'b110101000000?????????????1010011;
  localparam logic [31:0] FCVT_H_WU          = 32'b110101000001?????????????1010011;
  localparam logic [31:0] FMV_X_H            = 32'b111001000000?????000?????1010011;
  localparam logic [31:0] FCLASS_H           = 32'b111001000000?????001?????1010011;
  localparam logic [31:0] FMV_H_X            = 32'b111101000000?????000?????1010011;
  localparam logic [31:0] FCVT_L_H           = 32'b110001000010?????????????1010011;
  localparam logic [31:0] FCVT_LU_H          = 32'b110001000011?????????????1010011;
  localparam logic [31:0] FCVT_H_L           = 32'b110101000010?????????????1010011;
  localparam logic [31:0] FCVT_H_LU          = 32'b110101000011?????????????1010011;
  localparam logic [31:0] FCVT_S_H           = 32'b010000000010?????000?????1010011;
  localparam logic [31:0] FCVT_H_S           = 32'b010001000000?????????????1010011;
  localparam logic [31:0] FCVT_D_H           = 32'b010000100010?????000?????1010011;
  localparam logic [31:0] FCVT_H_D           = 32'b010001000001?????????????1010011;
  localparam logic [31:0] FLAH               = 32'b?????????????????001?????0000111;
  localparam logic [31:0] FSAH               = 32'b?????????????????001?????0100111;
  localparam logic [31:0] FMADD_AH           = 32'b?????10??????????????????1000011;
  localparam logic [31:0] FMSUB_AH           = 32'b?????10??????????????????1000111;
  localparam logic [31:0] FNMSUB_AH          = 32'b?????10??????????????????1001011;
  localparam logic [31:0] FNMADD_AH          = 32'b?????10??????????????????1001111;
  localparam logic [31:0] FADD_AH            = 32'b0000010??????????????????1010011;
  localparam logic [31:0] FSUB_AH            = 32'b0000110??????????????????1010011;
  localparam logic [31:0] FMUL_AH            = 32'b0001010??????????????????1010011;
  localparam logic [31:0] FDIV_AH            = 32'b0001110??????????????????1010011;
  localparam logic [31:0] FSQRT_AH           = 32'b010111000000?????????????1010011;
  localparam logic [31:0] FSGNJ_AH           = 32'b0010010??????????000?????1010011;
  localparam logic [31:0] FSGNJN_AH          = 32'b0010010??????????001?????1010011;
  localparam logic [31:0] FSGNJX_AH          = 32'b0010010??????????010?????1010011;
  localparam logic [31:0] FMIN_AH            = 32'b0010110??????????000?????1010011;
  localparam logic [31:0] FMAX_AH            = 32'b0010110??????????001?????1010011;
  localparam logic [31:0] FEQ_AH             = 32'b1010010??????????010?????1010011;
  localparam logic [31:0] FLT_AH             = 32'b1010010??????????001?????1010011;
  localparam logic [31:0] FLE_AH             = 32'b1010010??????????000?????1010011;
  localparam logic [31:0] FCVT_W_AH          = 32'b110001000000?????????????1010011;
  localparam logic [31:0] FCVT_WU_AH         = 32'b110001000001?????????????1010011;
  localparam logic [31:0] FCVT_AH_W          = 32'b110101000000?????????????1010011;
  localparam logic [31:0] FCVT_AH_WU         = 32'b110101000001?????????????1010011;
  localparam logic [31:0] FMV_X_AH           = 32'b111001000000?????000?????1010011;
  localparam logic [31:0] FCLASS_AH          = 32'b111001000000?????001?????1010011;
  localparam logic [31:0] FMV_AH_X           = 32'b111101000000?????000?????1010011;
  localparam logic [31:0] FCVT_L_AH          = 32'b110001000010?????????????1010011;
  localparam logic [31:0] FCVT_LU_AH         = 32'b110001000011?????????????1010011;
  localparam logic [31:0] FCVT_AH_L          = 32'b110101000010?????????????1010011;
  localparam logic [31:0] FCVT_AH_LU         = 32'b110101000011?????????????1010011;
  localparam logic [31:0] FCVT_S_AH          = 32'b010000000010?????000?????1010011;
  localparam logic [31:0] FCVT_AH_S          = 32'b010001000000?????????????1010011;
  localparam logic [31:0] FCVT_D_AH          = 32'b010000100010?????000?????1010011;
  localparam logic [31:0] FCVT_AH_D          = 32'b010001000001?????????????1010011;
  localparam logic [31:0] FCVT_H_H           = 32'b010001000010?????????????1010011;
  localparam logic [31:0] FCVT_AH_H          = 32'b010001000010?????????????1010011;
  localparam logic [31:0] FCVT_H_AH          = 32'b010001000010?????????????1010011;
  localparam logic [31:0] FCVT_AH_AH         = 32'b010001000010?????????????1010011;
  localparam logic [31:0] FLB                = 32'b?????????????????000?????0000111;
  localparam logic [31:0] FSB                = 32'b?????????????????000?????0100111;
  localparam logic [31:0] FMADD_B            = 32'b?????11??????????????????1000011;
  localparam logic [31:0] FMSUB_B            = 32'b?????11??????????????????1000111;
  localparam logic [31:0] FNMSUB_B           = 32'b?????11??????????????????1001011;
  localparam logic [31:0] FNMADD_B           = 32'b?????11??????????????????1001111;
  localparam logic [31:0] FADD_B             = 32'b0000011??????????????????1010011;
  localparam logic [31:0] FSUB_B             = 32'b0000111??????????????????1010011;
  localparam logic [31:0] FMUL_B             = 32'b0001011??????????????????1010011;
  localparam logic [31:0] FDIV_B             = 32'b0001111??????????????????1010011;
  localparam logic [31:0] FSQRT_B            = 32'b010111100000?????????????1010011;
  localparam logic [31:0] FSGNJ_B            = 32'b0010011??????????000?????1010011;
  localparam logic [31:0] FSGNJN_B           = 32'b0010011??????????001?????1010011;
  localparam logic [31:0] FSGNJX_B           = 32'b0010011??????????010?????1010011;
  localparam logic [31:0] FMIN_B             = 32'b0010111??????????000?????1010011;
  localparam logic [31:0] FMAX_B             = 32'b0010111??????????001?????1010011;
  localparam logic [31:0] FEQ_B              = 32'b1010011??????????010?????1010011;
  localparam logic [31:0] FLT_B              = 32'b1010011??????????001?????1010011;
  localparam logic [31:0] FLE_B              = 32'b1010011??????????000?????1010011;
  localparam logic [31:0] FCVT_W_B           = 32'b110001100000?????????????1010011;
  localparam logic [31:0] FCVT_WU_B          = 32'b110001100001?????????????1010011;
  localparam logic [31:0] FCVT_B_W           = 32'b110101100000?????????????1010011;
  localparam logic [31:0] FCVT_B_WU          = 32'b110101100001?????????????1010011;
  localparam logic [31:0] FMV_X_B            = 32'b111001100000?????000?????1010011;
  localparam logic [31:0] FCLASS_B           = 32'b111001100000?????001?????1010011;
  localparam logic [31:0] FMV_B_X            = 32'b111101100000?????000?????1010011;
  localparam logic [31:0] FCVT_L_B           = 32'b110001100010?????????????1010011;
  localparam logic [31:0] FCVT_LU_B          = 32'b110001100011?????????????1010011;
  localparam logic [31:0] FCVT_B_L           = 32'b110101100010?????????????1010011;
  localparam logic [31:0] FCVT_B_LU          = 32'b110101100011?????????????1010011;
  localparam logic [31:0] FCVT_S_B           = 32'b010000000011?????000?????1010011;
  localparam logic [31:0] FCVT_B_S           = 32'b010001100000?????????????1010011;
  localparam logic [31:0] FCVT_D_B           = 32'b010000100011?????000?????1010011;
  localparam logic [31:0] FCVT_B_D           = 32'b010001100001?????????????1010011;
  localparam logic [31:0] FCVT_H_B           = 32'b010001000011?????000?????1010011;
  localparam logic [31:0] FCVT_B_H           = 32'b010001100010?????????????1010011;
  localparam logic [31:0] FCVT_AH_B          = 32'b010001000011?????000?????1010011;
  localparam logic [31:0] FCVT_B_AH          = 32'b010001100010?????????????1010011;
  localparam logic [31:0] FLAB               = 32'b?????????????????000?????0000111;
  localparam logic [31:0] FSAB               = 32'b?????????????????000?????0100111;
  localparam logic [31:0] FMADD_AB           = 32'b?????11??????????????????1000011;
  localparam logic [31:0] FMSUB_AB           = 32'b?????11??????????????????1000111;
  localparam logic [31:0] FNMSUB_AB          = 32'b?????11??????????????????1001011;
  localparam logic [31:0] FNMADD_AB          = 32'b?????11??????????????????1001111;
  localparam logic [31:0] FADD_AB            = 32'b0000011??????????????????1010011;
  localparam logic [31:0] FSUB_AB            = 32'b0000111??????????????????1010011;
  localparam logic [31:0] FMUL_AB            = 32'b0001011??????????????????1010011;
  localparam logic [31:0] FDIV_AB            = 32'b0001111??????????????????1010011;
  localparam logic [31:0] FSQRT_AB           = 32'b010111100000?????????????1010011;
  localparam logic [31:0] FSGNJ_AB           = 32'b0010011??????????000?????1010011;
  localparam logic [31:0] FSGNJN_AB          = 32'b0010011??????????001?????1010011;
  localparam logic [31:0] FSGNJX_AB          = 32'b0010011??????????010?????1010011;
  localparam logic [31:0] FMIN_AB            = 32'b0010111??????????000?????1010011;
  localparam logic [31:0] FMAX_AB            = 32'b0010111??????????001?????1010011;
  localparam logic [31:0] FEQ_AB             = 32'b1010011??????????010?????1010011;
  localparam logic [31:0] FLT_AB             = 32'b1010011??????????001?????1010011;
  localparam logic [31:0] FLE_AB             = 32'b1010011??????????000?????1010011;
  localparam logic [31:0] FCVT_W_AB          = 32'b110001100000?????????????1010011;
  localparam logic [31:0] FCVT_WU_AB         = 32'b110001100001?????????????1010011;
  localparam logic [31:0] FCVT_AB_W          = 32'b110101100000?????????????1010011;
  localparam logic [31:0] FCVT_AB_WU         = 32'b110101100001?????????????1010011;
  localparam logic [31:0] FMV_X_AB           = 32'b111001100000?????000?????1010011;
  localparam logic [31:0] FCLASS_AB          = 32'b111001100000?????001?????1010011;
  localparam logic [31:0] FMV_AB_X           = 32'b111101100000?????000?????1010011;
  localparam logic [31:0] FCVT_L_AB          = 32'b110001100010?????????????1010011;
  localparam logic [31:0] FCVT_LU_AB         = 32'b110001100011?????????????1010011;
  localparam logic [31:0] FCVT_AB_L          = 32'b110101100010?????????????1010011;
  localparam logic [31:0] FCVT_AB_LU         = 32'b110101100011?????????????1010011;
  localparam logic [31:0] FCVT_S_AB          = 32'b010000000011?????000?????1010011;
  localparam logic [31:0] FCVT_AB_S          = 32'b010001100000?????????????1010011;
  localparam logic [31:0] FCVT_D_AB          = 32'b010000100011?????000?????1010011;
  localparam logic [31:0] FCVT_AB_D          = 32'b010001100001?????????????1010011;
  localparam logic [31:0] FCVT_H_AB          = 32'b010001000011?????000?????1010011;
  localparam logic [31:0] FCVT_AB_H          = 32'b010001100010?????????????1010011;
  localparam logic [31:0] FCVT_AH_AB         = 32'b010001000011?????000?????1010011;
  localparam logic [31:0] FCVT_AB_AH         = 32'b010001100010?????????????1010011;
  localparam logic [31:0] FCVT_B_B           = 32'b010001100011?????000?????1010011;
  localparam logic [31:0] FCVT_AB_B          = 32'b010001100011?????000?????1010011;
  localparam logic [31:0] FCVT_B_AB          = 32'b010001100011?????000?????1010011;
  localparam logic [31:0] FCVT_AB_AB         = 32'b010001100011?????000?????1010011;
  localparam logic [31:0] VFADD_S            = 32'b1000001??????????000?????0110011;
  localparam logic [31:0] VFADD_R_S          = 32'b1000001??????????100?????0110011;
  localparam logic [31:0] VFSUB_S            = 32'b1000010??????????000?????0110011;
  localparam logic [31:0] VFSUB_R_S          = 32'b1000010??????????100?????0110011;
  localparam logic [31:0] VFMUL_S            = 32'b1000011??????????000?????0110011;
  localparam logic [31:0] VFMUL_R_S          = 32'b1000011??????????100?????0110011;
  localparam logic [31:0] VFDIV_S            = 32'b1000100??????????000?????0110011;
  localparam logic [31:0] VFDIV_R_S          = 32'b1000100??????????100?????0110011;
  localparam logic [31:0] VFMIN_S            = 32'b1000101??????????000?????0110011;
  localparam logic [31:0] VFMIN_R_S          = 32'b1000101??????????100?????0110011;
  localparam logic [31:0] VFMAX_S            = 32'b1000110??????????000?????0110011;
  localparam logic [31:0] VFMAX_R_S          = 32'b1000110??????????100?????0110011;
  localparam logic [31:0] VFSQRT_S           = 32'b100011100000?????000?????0110011;
  localparam logic [31:0] VFMAC_S            = 32'b1001000??????????000?????0110011;
  localparam logic [31:0] VFMAC_R_S          = 32'b1001000??????????100?????0110011;
  localparam logic [31:0] VFMRE_S            = 32'b1001001??????????000?????0110011;
  localparam logic [31:0] VFMRE_R_S          = 32'b1001001??????????100?????0110011;
  localparam logic [31:0] VFCLASS_S          = 32'b100110000001?????000?????0110011;
  localparam logic [31:0] VFSGNJ_S           = 32'b1001101??????????000?????0110011;
  localparam logic [31:0] VFSGNJ_R_S         = 32'b1001101??????????100?????0110011;
  localparam logic [31:0] VFSGNJN_S          = 32'b1001110??????????000?????0110011;
  localparam logic [31:0] VFSGNJN_R_S        = 32'b1001110??????????100?????0110011;
  localparam logic [31:0] VFSGNJX_S          = 32'b1001111??????????000?????0110011;
  localparam logic [31:0] VFSGNJX_R_S        = 32'b1001111??????????100?????0110011;
  localparam logic [31:0] VFEQ_S             = 32'b1010000??????????000?????0110011;
  localparam logic [31:0] VFEQ_R_S           = 32'b1010000??????????100?????0110011;
  localparam logic [31:0] VFNE_S             = 32'b1010001??????????000?????0110011;
  localparam logic [31:0] VFNE_R_S           = 32'b1010001??????????100?????0110011;
  localparam logic [31:0] VFLT_S             = 32'b1010010??????????000?????0110011;
  localparam logic [31:0] VFLT_R_S           = 32'b1010010??????????100?????0110011;
  localparam logic [31:0] VFGE_S             = 32'b1010011??????????000?????0110011;
  localparam logic [31:0] VFGE_R_S           = 32'b1010011??????????100?????0110011;
  localparam logic [31:0] VFLE_S             = 32'b1010100??????????000?????0110011;
  localparam logic [31:0] VFLE_R_S           = 32'b1010100??????????100?????0110011;
  localparam logic [31:0] VFGT_S             = 32'b1010101??????????000?????0110011;
  localparam logic [31:0] VFGT_R_S           = 32'b1010101??????????100?????0110011;
  localparam logic [31:0] VFMV_X_S           = 32'b100110000000?????000?????0110011;
  localparam logic [31:0] VFMV_S_X           = 32'b100110000000?????100?????0110011;
  localparam logic [31:0] VFCVT_X_S          = 32'b100110000010?????000?????0110011;
  localparam logic [31:0] VFCVT_XU_S         = 32'b100110000010?????100?????0110011;
  localparam logic [31:0] VFCVT_S_X          = 32'b100110000011?????000?????0110011;
  localparam logic [31:0] VFCVT_S_XU         = 32'b100110000011?????100?????0110011;
  localparam logic [31:0] VFCPKA_S_S         = 32'b1011000??????????000?????0110011;
  localparam logic [31:0] VFCPKB_S_S         = 32'b1011000??????????100?????0110011;
  localparam logic [31:0] VFCPKC_S_S         = 32'b1011001??????????000?????0110011;
  localparam logic [31:0] VFCPKD_S_S         = 32'b1011001??????????100?????0110011;
  localparam logic [31:0] VFCPKA_S_D         = 32'b1011010??????????000?????0110011;
  localparam logic [31:0] VFCPKB_S_D         = 32'b1011010??????????100?????0110011;
  localparam logic [31:0] VFCPKC_S_D         = 32'b1011011??????????000?????0110011;
  localparam logic [31:0] VFCPKD_S_D         = 32'b1011011??????????100?????0110011;
  localparam logic [31:0] VFCVT_H_H          = 32'b100110000101?????010?????0110011;
  localparam logic [31:0] VFCVT_H_AH         = 32'b100110000101?????010?????0110011;
  localparam logic [31:0] VFCVT_AH_H         = 32'b100110000101?????010?????0110011;
  localparam logic [31:0] VFCVTU_H_H         = 32'b100110000101?????110?????0110011;
  localparam logic [31:0] VFCVTU_H_AH        = 32'b100110000101?????110?????0110011;
  localparam logic [31:0] VFCVTU_AH_H        = 32'b100110000101?????110?????0110011;
  localparam logic [31:0] VFADD_H            = 32'b1000001??????????010?????0110011;
  localparam logic [31:0] VFADD_R_H          = 32'b1000001??????????110?????0110011;
  localparam logic [31:0] VFSUB_H            = 32'b1000010??????????010?????0110011;
  localparam logic [31:0] VFSUB_R_H          = 32'b1000010??????????110?????0110011;
  localparam logic [31:0] VFMUL_H            = 32'b1000011??????????010?????0110011;
  localparam logic [31:0] VFMUL_R_H          = 32'b1000011??????????110?????0110011;
  localparam logic [31:0] VFDIV_H            = 32'b1000100??????????010?????0110011;
  localparam logic [31:0] VFDIV_R_H          = 32'b1000100??????????110?????0110011;
  localparam logic [31:0] VFMIN_H            = 32'b1000101??????????010?????0110011;
  localparam logic [31:0] VFMIN_R_H          = 32'b1000101??????????110?????0110011;
  localparam logic [31:0] VFMAX_H            = 32'b1000110??????????010?????0110011;
  localparam logic [31:0] VFMAX_R_H          = 32'b1000110??????????110?????0110011;
  localparam logic [31:0] VFSQRT_H           = 32'b100011100000?????010?????0110011;
  localparam logic [31:0] VFMAC_H            = 32'b1001000??????????010?????0110011;
  localparam logic [31:0] VFMAC_R_H          = 32'b1001000??????????110?????0110011;
  localparam logic [31:0] VFMRE_H            = 32'b1001001??????????010?????0110011;
  localparam logic [31:0] VFMRE_R_H          = 32'b1001001??????????110?????0110011;
  localparam logic [31:0] VFCLASS_H          = 32'b100110000001?????010?????0110011;
  localparam logic [31:0] VFSGNJ_H           = 32'b1001101??????????010?????0110011;
  localparam logic [31:0] VFSGNJ_R_H         = 32'b1001101??????????110?????0110011;
  localparam logic [31:0] VFSGNJN_H          = 32'b1001110??????????010?????0110011;
  localparam logic [31:0] VFSGNJN_R_H        = 32'b1001110??????????110?????0110011;
  localparam logic [31:0] VFSGNJX_H          = 32'b1001111??????????010?????0110011;
  localparam logic [31:0] VFSGNJX_R_H        = 32'b1001111??????????110?????0110011;
  localparam logic [31:0] VFEQ_H             = 32'b1010000??????????010?????0110011;
  localparam logic [31:0] VFEQ_R_H           = 32'b1010000??????????110?????0110011;
  localparam logic [31:0] VFNE_H             = 32'b1010001??????????010?????0110011;
  localparam logic [31:0] VFNE_R_H           = 32'b1010001??????????110?????0110011;
  localparam logic [31:0] VFLT_H             = 32'b1010010??????????010?????0110011;
  localparam logic [31:0] VFLT_R_H           = 32'b1010010??????????110?????0110011;
  localparam logic [31:0] VFGE_H             = 32'b1010011??????????010?????0110011;
  localparam logic [31:0] VFGE_R_H           = 32'b1010011??????????110?????0110011;
  localparam logic [31:0] VFLE_H             = 32'b1010100??????????010?????0110011;
  localparam logic [31:0] VFLE_R_H           = 32'b1010100??????????110?????0110011;
  localparam logic [31:0] VFGT_H             = 32'b1010101??????????010?????0110011;
  localparam logic [31:0] VFGT_R_H           = 32'b1010101??????????110?????0110011;
  localparam logic [31:0] VFMV_X_H           = 32'b100110000000?????010?????0110011;
  localparam logic [31:0] VFMV_H_X           = 32'b100110000000?????110?????0110011;
  localparam logic [31:0] VFCVT_X_H          = 32'b100110000010?????010?????0110011;
  localparam logic [31:0] VFCVT_XU_H         = 32'b100110000010?????110?????0110011;
  localparam logic [31:0] VFCVT_H_X          = 32'b100110000011?????010?????0110011;
  localparam logic [31:0] VFCVT_H_XU         = 32'b100110000011?????110?????0110011;
  localparam logic [31:0] VFCPKA_H_S         = 32'b1011000??????????010?????0110011;
  localparam logic [31:0] VFCPKB_H_S         = 32'b1011000??????????110?????0110011;
  localparam logic [31:0] VFCPKC_H_S         = 32'b1011001??????????010?????0110011;
  localparam logic [31:0] VFCPKD_H_S         = 32'b1011001??????????110?????0110011;
  localparam logic [31:0] VFCPKA_H_D         = 32'b1011010??????????010?????0110011;
  localparam logic [31:0] VFCPKB_H_D         = 32'b1011010??????????110?????0110011;
  localparam logic [31:0] VFCPKC_H_D         = 32'b1011011??????????010?????0110011;
  localparam logic [31:0] VFCPKD_H_D         = 32'b1011011??????????110?????0110011;
  localparam logic [31:0] VFCVT_S_H          = 32'b100110000110?????000?????0110011;
  localparam logic [31:0] VFCVTU_S_H         = 32'b100110000110?????100?????0110011;
  localparam logic [31:0] VFCVT_H_S          = 32'b100110000100?????010?????0110011;
  localparam logic [31:0] VFCVTU_H_S         = 32'b100110000100?????110?????0110011;
  localparam logic [31:0] VFADD_AH           = 32'b1000001??????????010?????0110011;
  localparam logic [31:0] VFADD_R_AH         = 32'b1000001??????????110?????0110011;
  localparam logic [31:0] VFSUB_AH           = 32'b1000010??????????010?????0110011;
  localparam logic [31:0] VFSUB_R_AH         = 32'b1000010??????????110?????0110011;
  localparam logic [31:0] VFMUL_AH           = 32'b1000011??????????010?????0110011;
  localparam logic [31:0] VFMUL_R_AH         = 32'b1000011??????????110?????0110011;
  localparam logic [31:0] VFDIV_AH           = 32'b1000100??????????010?????0110011;
  localparam logic [31:0] VFDIV_R_AH         = 32'b1000100??????????110?????0110011;
  localparam logic [31:0] VFMIN_AH           = 32'b1000101??????????010?????0110011;
  localparam logic [31:0] VFMIN_R_AH         = 32'b1000101??????????110?????0110011;
  localparam logic [31:0] VFMAX_AH           = 32'b1000110??????????010?????0110011;
  localparam logic [31:0] VFMAX_R_AH         = 32'b1000110??????????110?????0110011;
  localparam logic [31:0] VFSQRT_AH          = 32'b100011100000?????010?????0110011;
  localparam logic [31:0] VFMAC_AH           = 32'b1001000??????????010?????0110011;
  localparam logic [31:0] VFMAC_R_AH         = 32'b1001000??????????110?????0110011;
  localparam logic [31:0] VFMRE_AH           = 32'b1001001??????????010?????0110011;
  localparam logic [31:0] VFMRE_R_AH         = 32'b1001001??????????110?????0110011;
  localparam logic [31:0] VFCLASS_AH         = 32'b100110000001?????010?????0110011;
  localparam logic [31:0] VFSGNJ_AH          = 32'b1001101??????????010?????0110011;
  localparam logic [31:0] VFSGNJ_R_AH        = 32'b1001101??????????110?????0110011;
  localparam logic [31:0] VFSGNJN_AH         = 32'b1001110??????????010?????0110011;
  localparam logic [31:0] VFSGNJN_R_AH       = 32'b1001110??????????110?????0110011;
  localparam logic [31:0] VFSGNJX_AH         = 32'b1001111??????????010?????0110011;
  localparam logic [31:0] VFSGNJX_R_AH       = 32'b1001111??????????110?????0110011;
  localparam logic [31:0] VFEQ_AH            = 32'b1010000??????????010?????0110011;
  localparam logic [31:0] VFEQ_R_AH          = 32'b1010000??????????110?????0110011;
  localparam logic [31:0] VFNE_AH            = 32'b1010001??????????010?????0110011;
  localparam logic [31:0] VFNE_R_AH          = 32'b1010001??????????110?????0110011;
  localparam logic [31:0] VFLT_AH            = 32'b1010010??????????010?????0110011;
  localparam logic [31:0] VFLT_R_AH          = 32'b1010010??????????110?????0110011;
  localparam logic [31:0] VFGE_AH            = 32'b1010011??????????010?????0110011;
  localparam logic [31:0] VFGE_R_AH          = 32'b1010011??????????110?????0110011;
  localparam logic [31:0] VFLE_AH            = 32'b1010100??????????010?????0110011;
  localparam logic [31:0] VFLE_R_AH          = 32'b1010100??????????110?????0110011;
  localparam logic [31:0] VFGT_AH            = 32'b1010101??????????010?????0110011;
  localparam logic [31:0] VFGT_R_AH          = 32'b1010101??????????110?????0110011;
  localparam logic [31:0] VFMV_X_AH          = 32'b100110000000?????010?????0110011;
  localparam logic [31:0] VFMV_AH_X          = 32'b100110000000?????110?????0110011;
  localparam logic [31:0] VFCVT_X_AH         = 32'b100110000010?????010?????0110011;
  localparam logic [31:0] VFCVT_XU_AH        = 32'b100110000010?????110?????0110011;
  localparam logic [31:0] VFCVT_AH_X         = 32'b100110000011?????010?????0110011;
  localparam logic [31:0] VFCVT_AH_XU        = 32'b100110000011?????110?????0110011;
  localparam logic [31:0] VFCPKA_AH_S        = 32'b1011000??????????010?????0110011;
  localparam logic [31:0] VFCPKB_AH_S        = 32'b1011000??????????110?????0110011;
  localparam logic [31:0] VFCPKC_AH_S        = 32'b1011001??????????010?????0110011;
  localparam logic [31:0] VFCPKD_AH_S        = 32'b1011001??????????110?????0110011;
  localparam logic [31:0] VFCPKA_AH_D        = 32'b1011010??????????010?????0110011;
  localparam logic [31:0] VFCPKB_AH_D        = 32'b1011010??????????110?????0110011;
  localparam logic [31:0] VFCPKC_AH_D        = 32'b1011011??????????010?????0110011;
  localparam logic [31:0] VFCPKD_AH_D        = 32'b1011011??????????110?????0110011;
  localparam logic [31:0] VFCVT_S_AH         = 32'b100110000110?????000?????0110011;
  localparam logic [31:0] VFCVTU_S_AH        = 32'b100110000110?????100?????0110011;
  localparam logic [31:0] VFCVT_AH_S         = 32'b100110000100?????010?????0110011;
  localparam logic [31:0] VFCVTU_AH_S        = 32'b100110000100?????110?????0110011;
  localparam logic [31:0] VFADD_B            = 32'b1000001??????????011?????0110011;
  localparam logic [31:0] VFADD_R_B          = 32'b1000001??????????111?????0110011;
  localparam logic [31:0] VFSUB_B            = 32'b1000010??????????011?????0110011;
  localparam logic [31:0] VFSUB_R_B          = 32'b1000010??????????111?????0110011;
  localparam logic [31:0] VFMUL_B            = 32'b1000011??????????011?????0110011;
  localparam logic [31:0] VFMUL_R_B          = 32'b1000011??????????111?????0110011;
  localparam logic [31:0] VFDIV_B            = 32'b1000100??????????011?????0110011;
  localparam logic [31:0] VFDIV_R_B          = 32'b1000100??????????111?????0110011;
  localparam logic [31:0] VFMIN_B            = 32'b1000101??????????011?????0110011;
  localparam logic [31:0] VFMIN_R_B          = 32'b1000101??????????111?????0110011;
  localparam logic [31:0] VFMAX_B            = 32'b1000110??????????011?????0110011;
  localparam logic [31:0] VFMAX_R_B          = 32'b1000110??????????111?????0110011;
  localparam logic [31:0] VFSQRT_B           = 32'b100011100000?????011?????0110011;
  localparam logic [31:0] VFMAC_B            = 32'b1001000??????????011?????0110011;
  localparam logic [31:0] VFMAC_R_B          = 32'b1001000??????????111?????0110011;
  localparam logic [31:0] VFMRE_B            = 32'b1001001??????????011?????0110011;
  localparam logic [31:0] VFMRE_R_B          = 32'b1001001??????????111?????0110011;
  localparam logic [31:0] VFSGNJ_B           = 32'b1001101??????????011?????0110011;
  localparam logic [31:0] VFSGNJ_R_B         = 32'b1001101??????????111?????0110011;
  localparam logic [31:0] VFSGNJN_B          = 32'b1001110??????????011?????0110011;
  localparam logic [31:0] VFSGNJN_R_B        = 32'b1001110??????????111?????0110011;
  localparam logic [31:0] VFSGNJX_B          = 32'b1001111??????????011?????0110011;
  localparam logic [31:0] VFSGNJX_R_B        = 32'b1001111??????????111?????0110011;
  localparam logic [31:0] VFEQ_B             = 32'b1010000??????????011?????0110011;
  localparam logic [31:0] VFEQ_R_B           = 32'b1010000??????????111?????0110011;
  localparam logic [31:0] VFNE_B             = 32'b1010001??????????011?????0110011;
  localparam logic [31:0] VFNE_R_B           = 32'b1010001??????????111?????0110011;
  localparam logic [31:0] VFLT_B             = 32'b1010010??????????011?????0110011;
  localparam logic [31:0] VFLT_R_B           = 32'b1010010??????????111?????0110011;
  localparam logic [31:0] VFGE_B             = 32'b1010011??????????011?????0110011;
  localparam logic [31:0] VFGE_R_B           = 32'b1010011??????????111?????0110011;
  localparam logic [31:0] VFLE_B             = 32'b1010100??????????011?????0110011;
  localparam logic [31:0] VFLE_R_B           = 32'b1010100??????????111?????0110011;
  localparam logic [31:0] VFGT_B             = 32'b1010101??????????011?????0110011;
  localparam logic [31:0] VFGT_R_B           = 32'b1010101??????????111?????0110011;
  localparam logic [31:0] VFMV_X_B           = 32'b100110000000?????011?????0110011;
  localparam logic [31:0] VFMV_B_X           = 32'b100110000000?????111?????0110011;
  localparam logic [31:0] VFCLASS_B          = 32'b100110000001?????011?????0110011;
  localparam logic [31:0] VFCVT_X_B          = 32'b100110000010?????011?????0110011;
  localparam logic [31:0] VFCVT_XU_B         = 32'b100110000010?????111?????0110011;
  localparam logic [31:0] VFCVT_B_X          = 32'b100110000011?????011?????0110011;
  localparam logic [31:0] VFCVT_B_XU         = 32'b100110000011?????111?????0110011;
  localparam logic [31:0] VFCPKA_B_S         = 32'b1011000??????????011?????0110011;
  localparam logic [31:0] VFCPKB_B_S         = 32'b1011000??????????111?????0110011;
  localparam logic [31:0] VFCPKC_B_S         = 32'b1011001??????????011?????0110011;
  localparam logic [31:0] VFCPKD_B_S         = 32'b1011001??????????111?????0110011;
  localparam logic [31:0] VFCPKA_B_D         = 32'b1011010??????????011?????0110011;
  localparam logic [31:0] VFCPKB_B_D         = 32'b1011010??????????111?????0110011;
  localparam logic [31:0] VFCPKC_B_D         = 32'b1011011??????????011?????0110011;
  localparam logic [31:0] VFCPKD_B_D         = 32'b1011011??????????111?????0110011;
  localparam logic [31:0] VFCVT_S_B          = 32'b100110000111?????000?????0110011;
  localparam logic [31:0] VFCVTU_S_B         = 32'b100110000111?????100?????0110011;
  localparam logic [31:0] VFCVT_B_S          = 32'b100110000100?????011?????0110011;
  localparam logic [31:0] VFCVTU_B_S         = 32'b100110000100?????111?????0110011;
  localparam logic [31:0] VFCVT_H_B          = 32'b100110000111?????010?????0110011;
  localparam logic [31:0] VFCVTU_H_B         = 32'b100110000111?????110?????0110011;
  localparam logic [31:0] VFCVT_B_H          = 32'b100110000110?????011?????0110011;
  localparam logic [31:0] VFCVTU_B_H         = 32'b100110000110?????111?????0110011;
  localparam logic [31:0] VFCVT_AH_B         = 32'b100110000111?????010?????0110011;
  localparam logic [31:0] VFCVTU_AH_B        = 32'b100110000111?????110?????0110011;
  localparam logic [31:0] VFCVT_B_AH         = 32'b100110000110?????011?????0110011;
  localparam logic [31:0] VFCVTU_B_AH        = 32'b100110000110?????111?????0110011;
  localparam logic [31:0] VFCVT_B_B          = 32'b100110000111?????011?????0110011;
  localparam logic [31:0] VFCVT_AB_B         = 32'b100110000111?????011?????0110011;
  localparam logic [31:0] VFCVT_B_AB         = 32'b100110000111?????011?????0110011;
  localparam logic [31:0] VFCVTU_B_B         = 32'b100110000111?????111?????0110011;
  localparam logic [31:0] VFCVTU_AB_B        = 32'b100110000111?????111?????0110011;
  localparam logic [31:0] VFCVTU_B_AB        = 32'b100110000111?????111?????0110011;
  localparam logic [31:0] VFADD_AB           = 32'b1000001??????????011?????0110011;
  localparam logic [31:0] VFADD_R_AB         = 32'b1000001??????????111?????0110011;
  localparam logic [31:0] VFSUB_AB           = 32'b1000010??????????011?????0110011;
  localparam logic [31:0] VFSUB_R_AB         = 32'b1000010??????????111?????0110011;
  localparam logic [31:0] VFMUL_AB           = 32'b1000011??????????011?????0110011;
  localparam logic [31:0] VFMUL_R_AB         = 32'b1000011??????????111?????0110011;
  localparam logic [31:0] VFDIV_AB           = 32'b1000100??????????011?????0110011;
  localparam logic [31:0] VFDIV_R_AB         = 32'b1000100??????????111?????0110011;
  localparam logic [31:0] VFMIN_AB           = 32'b1000101??????????011?????0110011;
  localparam logic [31:0] VFMIN_R_AB         = 32'b1000101??????????111?????0110011;
  localparam logic [31:0] VFMAX_AB           = 32'b1000110??????????011?????0110011;
  localparam logic [31:0] VFMAX_R_AB         = 32'b1000110??????????111?????0110011;
  localparam logic [31:0] VFSQRT_AB          = 32'b100011100000?????011?????0110011;
  localparam logic [31:0] VFMAC_AB           = 32'b1001000??????????011?????0110011;
  localparam logic [31:0] VFMAC_R_AB         = 32'b1001000??????????111?????0110011;
  localparam logic [31:0] VFMRE_AB           = 32'b1001001??????????011?????0110011;
  localparam logic [31:0] VFMRE_R_AB         = 32'b1001001??????????111?????0110011;
  localparam logic [31:0] VFSGNJ_AB          = 32'b1001101??????????011?????0110011;
  localparam logic [31:0] VFSGNJ_R_AB        = 32'b1001101??????????111?????0110011;
  localparam logic [31:0] VFSGNJN_AB         = 32'b1001110??????????011?????0110011;
  localparam logic [31:0] VFSGNJN_R_AB       = 32'b1001110??????????111?????0110011;
  localparam logic [31:0] VFSGNJX_AB         = 32'b1001111??????????011?????0110011;
  localparam logic [31:0] VFSGNJX_R_AB       = 32'b1001111??????????111?????0110011;
  localparam logic [31:0] VFEQ_AB            = 32'b1010000??????????011?????0110011;
  localparam logic [31:0] VFEQ_R_AB          = 32'b1010000??????????111?????0110011;
  localparam logic [31:0] VFNE_AB            = 32'b1010001??????????011?????0110011;
  localparam logic [31:0] VFNE_R_AB          = 32'b1010001??????????111?????0110011;
  localparam logic [31:0] VFLT_AB            = 32'b1010010??????????011?????0110011;
  localparam logic [31:0] VFLT_R_AB          = 32'b1010010??????????111?????0110011;
  localparam logic [31:0] VFGE_AB            = 32'b1010011??????????011?????0110011;
  localparam logic [31:0] VFGE_R_AB          = 32'b1010011??????????111?????0110011;
  localparam logic [31:0] VFLE_AB            = 32'b1010100??????????011?????0110011;
  localparam logic [31:0] VFLE_R_AB          = 32'b1010100??????????111?????0110011;
  localparam logic [31:0] VFGT_AB            = 32'b1010101??????????011?????0110011;
  localparam logic [31:0] VFGT_R_AB          = 32'b1010101??????????111?????0110011;
  localparam logic [31:0] VFMV_X_AB          = 32'b100110000000?????011?????0110011;
  localparam logic [31:0] VFMV_AB_X          = 32'b100110000000?????111?????0110011;
  localparam logic [31:0] VFCLASS_AB         = 32'b100110000001?????011?????0110011;
  localparam logic [31:0] VFCVT_X_AB         = 32'b100110000010?????011?????0110011;
  localparam logic [31:0] VFCVT_XU_AB        = 32'b100110000010?????111?????0110011;
  localparam logic [31:0] VFCVT_AB_X         = 32'b100110000011?????011?????0110011;
  localparam logic [31:0] VFCVT_AB_XU        = 32'b100110000011?????111?????0110011;
  localparam logic [31:0] VFCPKA_AB_S        = 32'b1011000??????????011?????0110011;
  localparam logic [31:0] VFCPKB_AB_S        = 32'b1011000??????????111?????0110011;
  localparam logic [31:0] VFCPKC_AB_S        = 32'b1011001??????????011?????0110011;
  localparam logic [31:0] VFCPKD_AB_S        = 32'b1011001??????????111?????0110011;
  localparam logic [31:0] VFCPKA_AB_D        = 32'b1011010??????????011?????0110011;
  localparam logic [31:0] VFCPKB_AB_D        = 32'b1011010??????????111?????0110011;
  localparam logic [31:0] VFCPKC_AB_D        = 32'b1011011??????????011?????0110011;
  localparam logic [31:0] VFCPKD_AB_D        = 32'b1011011??????????111?????0110011;
  localparam logic [31:0] VFCVT_S_AB         = 32'b100110000111?????000?????0110011;
  localparam logic [31:0] VFCVTU_S_AB        = 32'b100110000111?????100?????0110011;
  localparam logic [31:0] VFCVT_AB_S         = 32'b100110000100?????011?????0110011;
  localparam logic [31:0] VFCVTU_AB_S        = 32'b100110000100?????111?????0110011;
  localparam logic [31:0] VFCVT_H_AB         = 32'b100110000111?????010?????0110011;
  localparam logic [31:0] VFCVTU_H_AB        = 32'b100110000111?????110?????0110011;
  localparam logic [31:0] VFCVT_AB_H         = 32'b100110000110?????011?????0110011;
  localparam logic [31:0] VFCVTU_AB_H        = 32'b100110000110?????111?????0110011;
  localparam logic [31:0] VFCVT_AH_AB        = 32'b100110000111?????010?????0110011;
  localparam logic [31:0] VFCVTU_AH_AB       = 32'b100110000111?????110?????0110011;
  localparam logic [31:0] VFCVT_AB_AH        = 32'b100110000110?????011?????0110011;
  localparam logic [31:0] VFCVTU_AB_AH       = 32'b100110000110?????111?????0110011;
  localparam logic [31:0] FMULEX_S_H         = 32'b0100110??????????????????1010011;
  localparam logic [31:0] FMACEX_S_H         = 32'b0101010??????????????????1010011;
  localparam logic [31:0] FMULEX_S_AH        = 32'b0100110??????????????????1010011;
  localparam logic [31:0] FMACEX_S_AH        = 32'b0101010??????????????????1010011;
  localparam logic [31:0] FMULEX_S_B         = 32'b0100111??????????????????1010011;
  localparam logic [31:0] FMACEX_S_B         = 32'b0101011??????????????????1010011;
  localparam logic [31:0] FMULEX_S_AB        = 32'b0100111??????????????????1010011;
  localparam logic [31:0] FMACEX_S_AB        = 32'b0101011??????????????????1010011;
  localparam logic [31:0] VFSUM_S            = 32'b100011111100?????000?????0110011;
  localparam logic [31:0] VFNSUM_S           = 32'b101011111100?????000?????0110011;
  localparam logic [31:0] VFSUM_H            = 32'b100011111110?????010?????0110011;
  localparam logic [31:0] VFNSUM_H           = 32'b101011111110?????010?????0110011;
  localparam logic [31:0] VFSUM_AH           = 32'b100011111110?????010?????0110011;
  localparam logic [31:0] VFNSUM_AH          = 32'b101011111110?????010?????0110011;
  localparam logic [31:0] VFSUM_B            = 32'b100011100111?????011?????0110011;
  localparam logic [31:0] VFNSUM_B           = 32'b101011100111?????011?????0110011;
  localparam logic [31:0] VFSUM_AB           = 32'b100011100111?????011?????0110011;
  localparam logic [31:0] VFNSUM_AB          = 32'b101011100111?????011?????0110011;
  localparam logic [31:0] VFSUMEX_S_H        = 32'b100011110110?????000?????0110011;
  localparam logic [31:0] VFNSUMEX_S_H       = 32'b101011110110?????000?????0110011;
  localparam logic [31:0] VFDOTPEX_S_H       = 32'b1001011??????????000?????0110011;
  localparam logic [31:0] VFDOTPEX_S_R_H     = 32'b1001011??????????100?????0110011;
  localparam logic [31:0] VFNDOTPEX_S_H      = 32'b1011101??????????000?????0110011;
  localparam logic [31:0] VFNDOTPEX_S_R_H    = 32'b1011101??????????100?????0110011;
  localparam logic [31:0] VFSUMEX_S_AH       = 32'b100011110110?????000?????0110011;
  localparam logic [31:0] VFNSUMEX_S_AH      = 32'b101011110110?????000?????0110011;
  localparam logic [31:0] VFDOTPEX_S_AH      = 32'b1001011??????????000?????0110011;
  localparam logic [31:0] VFDOTPEX_S_R_AH    = 32'b1001011??????????100?????0110011;
  localparam logic [31:0] VFNDOTPEX_S_AH     = 32'b1011101??????????000?????0110011;
  localparam logic [31:0] VFNDOTPEX_S_R_AH   = 32'b1011101??????????100?????0110011;
  localparam logic [31:0] VFSUMEX_H_B        = 32'b100011110111?????010?????0110011;
  localparam logic [31:0] VFNSUMEX_H_B       = 32'b101011110111?????010?????0110011;
  localparam logic [31:0] VFDOTPEX_H_B       = 32'b1001011??????????010?????0110011;
  localparam logic [31:0] VFDOTPEX_H_R_B     = 32'b1001011??????????110?????0110011;
  localparam logic [31:0] VFNDOTPEX_H_B      = 32'b1011101??????????010?????0110011;
  localparam logic [31:0] VFNDOTPEX_H_R_B    = 32'b1011101??????????110?????0110011;
  localparam logic [31:0] VFSUMEX_AH_B       = 32'b100011110111?????010?????0110011;
  localparam logic [31:0] VFNSUMEX_AH_B      = 32'b101011110111?????010?????0110011;
  localparam logic [31:0] VFDOTPEX_AH_B      = 32'b1001011??????????010?????0110011;
  localparam logic [31:0] VFDOTPEX_AH_R_B    = 32'b1001011??????????110?????0110011;
  localparam logic [31:0] VFNDOTPEX_AH_B     = 32'b1011101??????????010?????0110011;
  localparam logic [31:0] VFNDOTPEX_AH_R_B   = 32'b1011101??????????110?????0110011;
  localparam logic [31:0] VFSUMEX_H_AB       = 32'b100011110111?????010?????0110011;
  localparam logic [31:0] VFNSUMEX_H_AB      = 32'b101011110111?????010?????0110011;
  localparam logic [31:0] VFDOTPEX_H_AB      = 32'b1001011??????????010?????0110011;
  localparam logic [31:0] VFDOTPEX_H_R_AB    = 32'b1001011??????????110?????0110011;
  localparam logic [31:0] VFNDOTPEX_H_AB     = 32'b1011101??????????010?????0110011;
  localparam logic [31:0] VFNDOTPEX_H_R_AB   = 32'b1011101??????????110?????0110011;
  localparam logic [31:0] VFSUMEX_AH_AB      = 32'b100011110111?????010?????0110011;
  localparam logic [31:0] VFNSUMEX_AH_AB     = 32'b101011110111?????010?????0110011;
  localparam logic [31:0] VFDOTPEX_AH_AB     = 32'b1001011??????????010?????0110011;
  localparam logic [31:0] VFDOTPEX_AH_R_AB   = 32'b1001011??????????110?????0110011;
  localparam logic [31:0] VFNDOTPEX_AH_AB    = 32'b1011101??????????010?????0110011;
  localparam logic [31:0] VFNDOTPEX_AH_R_AB  = 32'b1011101??????????110?????0110011;
  localparam logic [31:0] IMV_X_W            = 32'b111000000000?????000?????1011011;
  localparam logic [31:0] IMV_W_X            = 32'b111100000000?????000?????1011011;
  localparam logic [31:0] IADDI              = 32'b?????????????????000?????1111011;
  localparam logic [31:0] ISLLI              = 32'b000000???????????001?????1111011;
  localparam logic [31:0] ISLTI              = 32'b?????????????????010?????1111011;
  localparam logic [31:0] ISLTIU             = 32'b?????????????????011?????1111011;
  localparam logic [31:0] IXORI              = 32'b?????????????????100?????1111011;
  localparam logic [31:0] ISRLI              = 32'b000000???????????101?????1111011;
  localparam logic [31:0] ISRAI              = 32'b010000???????????101?????1111011;
  localparam logic [31:0] IORI               = 32'b?????????????????110?????1111011;
  localparam logic [31:0] IANDI              = 32'b?????????????????111?????1111011;
  localparam logic [31:0] IADD               = 32'b0000000??????????000?????1011011;
  localparam logic [31:0] ISUB               = 32'b0100000??????????000?????1011011;
  localparam logic [31:0] ISLL               = 32'b0000000??????????001?????1011011;
  localparam logic [31:0] ISLT               = 32'b0000000??????????010?????1011011;
  localparam logic [31:0] ISLTU              = 32'b0000000??????????011?????1011011;
  localparam logic [31:0] IXOR               = 32'b0000000??????????100?????1011011;
  localparam logic [31:0] ISRL               = 32'b0000000??????????101?????1011011;
  localparam logic [31:0] ISRA               = 32'b0100000??????????101?????1011011;
  localparam logic [31:0] IOR                = 32'b0000000??????????110?????1011011;
  localparam logic [31:0] IAND               = 32'b0000000??????????111?????1011011;
  localparam logic [31:0] IMADD              = 32'b?????01??????????000?????1011011;
  localparam logic [31:0] IMSUB              = 32'b?????01??????????001?????1011011;
  localparam logic [31:0] INMSUB             = 32'b?????01??????????010?????1011011;
  localparam logic [31:0] INMADD             = 32'b?????01??????????011?????1011011;
  localparam logic [31:0] IMUL               = 32'b0000010??????????000?????1011011;
  localparam logic [31:0] IMULH              = 32'b0000010??????????001?????1011011;
  localparam logic [31:0] IMULHSU            = 32'b0000010??????????010?????1011011;
  localparam logic [31:0] IMULHU             = 32'b0000010??????????011?????1011011;
  localparam logic [31:0] IANDN              = 32'b0100000??????????111?????1011011;
  localparam logic [31:0] IORN               = 32'b0100000??????????110?????1011011;
  localparam logic [31:0] IXNOR              = 32'b0100000??????????100?????1011011;
  localparam logic [31:0] ISLO               = 32'b0010000??????????001?????1011011;
  localparam logic [31:0] ISRO               = 32'b0010000??????????101?????1011011;
  localparam logic [31:0] IROL               = 32'b0110000??????????001?????1011011;
  localparam logic [31:0] IROR               = 32'b0110000??????????101?????1011011;
  localparam logic [31:0] ISBCLR             = 32'b0100100??????????001?????1011011;
  localparam logic [31:0] ISBSET             = 32'b0010100??????????001?????1011011;
  localparam logic [31:0] ISBINV             = 32'b0110100??????????001?????1011011;
  localparam logic [31:0] ISBEXT             = 32'b0100100??????????101?????1011011;
  localparam logic [31:0] IGORC              = 32'b0010100??????????101?????1011011;
  localparam logic [31:0] IGREV              = 32'b0110100??????????101?????1011011;
  localparam logic [31:0] ISLOI              = 32'b001000???????????001?????1111011;
  localparam logic [31:0] ISROI              = 32'b001000???????????101?????1111011;
  localparam logic [31:0] IRORI              = 32'b011000???????????101?????1111011;
  localparam logic [31:0] ISBCLRI            = 32'b010010???????????001?????1111011;
  localparam logic [31:0] ISBSETI            = 32'b001010???????????001?????1111011;
  localparam logic [31:0] ISBINVI            = 32'b011010???????????001?????1111011;
  localparam logic [31:0] ISBEXTI            = 32'b010010???????????101?????1111011;
  localparam logic [31:0] IGORCI             = 32'b001010???????????101?????1111011;
  localparam logic [31:0] IGREVI             = 32'b011010???????????101?????1111011;
  localparam logic [31:0] ICLZ               = 32'b011000000000?????010?????1011011;
  localparam logic [31:0] ICTZ               = 32'b011000000001?????010?????1011011;
  localparam logic [31:0] IPCNT              = 32'b011000000010?????010?????1011011;
  localparam logic [31:0] ISEXT_B            = 32'b011000000100?????010?????1011011;
  localparam logic [31:0] ISEXT_H            = 32'b011000000101?????010?????1011011;
  localparam logic [31:0] ICRC32_B           = 32'b011000010000?????001?????1011011;
  localparam logic [31:0] ICRC32_H           = 32'b011000010001?????001?????1011011;
  localparam logic [31:0] ICRC32_W           = 32'b011000010010?????001?????1011011;
  localparam logic [31:0] ICRC32C_B          = 32'b011000011000?????001?????1011011;
  localparam logic [31:0] ICRC32C_H          = 32'b011000011001?????001?????1011011;
  localparam logic [31:0] ICRC32C_W          = 32'b011000011010?????001?????1011011;
  localparam logic [31:0] ISH1ADD            = 32'b0010000??????????010?????1011011;
  localparam logic [31:0] ISH2ADD            = 32'b0010000??????????100?????1011011;
  localparam logic [31:0] ISH3ADD            = 32'b0010000??????????110?????1011011;
  localparam logic [31:0] ICLMUL             = 32'b0000101??????????001?????1011011;
  localparam logic [31:0] ICLMULR            = 32'b0000101??????????010?????1011011;
  localparam logic [31:0] ICLMULH            = 32'b0000101??????????011?????1011011;
  localparam logic [31:0] IMIN               = 32'b0000101??????????100?????1011011;
  localparam logic [31:0] IMAX               = 32'b0000101??????????101?????1011011;
  localparam logic [31:0] IMINU              = 32'b0000101??????????110?????1011011;
  localparam logic [31:0] IMAXU              = 32'b0000101??????????111?????1011011;
  localparam logic [31:0] ISHFL              = 32'b0000100??????????001?????1011011;
  localparam logic [31:0] IUNSHFL            = 32'b0000100??????????101?????1011011;
  localparam logic [31:0] IBEXT              = 32'b0000100??????????110?????1011011;
  localparam logic [31:0] IBDEP              = 32'b0100100??????????110?????1011011;
  localparam logic [31:0] IPACK              = 32'b0000100??????????100?????1011011;
  localparam logic [31:0] IPACKU             = 32'b0100100??????????100?????1011011;
  localparam logic [31:0] IPACKH             = 32'b0000100??????????111?????1011011;
  localparam logic [31:0] IBFP               = 32'b0100100??????????111?????1011011;
  localparam logic [31:0] ISHFLI             = 32'b0000100??????????001?????1111011;
  localparam logic [31:0] IUNSHFLI           = 32'b0000100??????????101?????1111011;
  /* CSR Addresses */
  localparam logic [11:0] CSR_FFLAGS = 12'h1;
  localparam logic [11:0] CSR_FRM = 12'h2;
  localparam logic [11:0] CSR_FCSR = 12'h3;
  localparam logic [11:0] CSR_FMODE = 12'h800;
  localparam logic [11:0] CSR_FSRM = 12'h801;
  localparam logic [11:0] CSR_CYCLE = 12'hc00;
  localparam logic [11:0] CSR_TIME = 12'hc01;
  localparam logic [11:0] CSR_INSTRET = 12'hc02;
  localparam logic [11:0] CSR_HPMCOUNTER3 = 12'hc03;
  localparam logic [11:0] CSR_HPMCOUNTER4 = 12'hc04;
  localparam logic [11:0] CSR_HPMCOUNTER5 = 12'hc05;
  localparam logic [11:0] CSR_HPMCOUNTER6 = 12'hc06;
  localparam logic [11:0] CSR_HPMCOUNTER7 = 12'hc07;
  localparam logic [11:0] CSR_HPMCOUNTER8 = 12'hc08;
  localparam logic [11:0] CSR_HPMCOUNTER9 = 12'hc09;
  localparam logic [11:0] CSR_HPMCOUNTER10 = 12'hc0a;
  localparam logic [11:0] CSR_HPMCOUNTER11 = 12'hc0b;
  localparam logic [11:0] CSR_HPMCOUNTER12 = 12'hc0c;
  localparam logic [11:0] CSR_HPMCOUNTER13 = 12'hc0d;
  localparam logic [11:0] CSR_HPMCOUNTER14 = 12'hc0e;
  localparam logic [11:0] CSR_HPMCOUNTER15 = 12'hc0f;
  localparam logic [11:0] CSR_HPMCOUNTER16 = 12'hc10;
  localparam logic [11:0] CSR_HPMCOUNTER17 = 12'hc11;
  localparam logic [11:0] CSR_HPMCOUNTER18 = 12'hc12;
  localparam logic [11:0] CSR_HPMCOUNTER19 = 12'hc13;
  localparam logic [11:0] CSR_HPMCOUNTER20 = 12'hc14;
  localparam logic [11:0] CSR_HPMCOUNTER21 = 12'hc15;
  localparam logic [11:0] CSR_HPMCOUNTER22 = 12'hc16;
  localparam logic [11:0] CSR_HPMCOUNTER23 = 12'hc17;
  localparam logic [11:0] CSR_HPMCOUNTER24 = 12'hc18;
  localparam logic [11:0] CSR_HPMCOUNTER25 = 12'hc19;
  localparam logic [11:0] CSR_HPMCOUNTER26 = 12'hc1a;
  localparam logic [11:0] CSR_HPMCOUNTER27 = 12'hc1b;
  localparam logic [11:0] CSR_HPMCOUNTER28 = 12'hc1c;
  localparam logic [11:0] CSR_HPMCOUNTER29 = 12'hc1d;
  localparam logic [11:0] CSR_HPMCOUNTER30 = 12'hc1e;
  localparam logic [11:0] CSR_HPMCOUNTER31 = 12'hc1f;
  localparam logic [11:0] CSR_SSTATUS = 12'h100;
  localparam logic [11:0] CSR_SIE = 12'h104;
  localparam logic [11:0] CSR_STVEC = 12'h105;
  localparam logic [11:0] CSR_SCOUNTEREN = 12'h106;
  localparam logic [11:0] CSR_SSCRATCH = 12'h140;
  localparam logic [11:0] CSR_SEPC = 12'h141;
  localparam logic [11:0] CSR_SCAUSE = 12'h142;
  localparam logic [11:0] CSR_STVAL = 12'h143;
  localparam logic [11:0] CSR_SIP = 12'h144;
  localparam logic [11:0] CSR_SATP = 12'h180;
  localparam logic [11:0] CSR_BSSTATUS = 12'h200;
  localparam logic [11:0] CSR_BSIE = 12'h204;
  localparam logic [11:0] CSR_BSTVEC = 12'h205;
  localparam logic [11:0] CSR_BSSCRATCH = 12'h240;
  localparam logic [11:0] CSR_BSEPC = 12'h241;
  localparam logic [11:0] CSR_BSCAUSE = 12'h242;
  localparam logic [11:0] CSR_BSTVAL = 12'h243;
  localparam logic [11:0] CSR_BSIP = 12'h244;
  localparam logic [11:0] CSR_BSATP = 12'h280;
  localparam logic [11:0] CSR_HSTATUS = 12'ha00;
  localparam logic [11:0] CSR_HEDELEG = 12'ha02;
  localparam logic [11:0] CSR_HIDELEG = 12'ha03;
  localparam logic [11:0] CSR_HGATP = 12'ha80;
  localparam logic [11:0] CSR_UTVT = 12'h7;
  localparam logic [11:0] CSR_UNXTI = 12'h45;
  localparam logic [11:0] CSR_UINTSTATUS = 12'h46;
  localparam logic [11:0] CSR_USCRATCHCSW = 12'h48;
  localparam logic [11:0] CSR_USCRATCHCSWL = 12'h49;
  localparam logic [11:0] CSR_STVT = 12'h107;
  localparam logic [11:0] CSR_SNXTI = 12'h145;
  localparam logic [11:0] CSR_SINTSTATUS = 12'h146;
  localparam logic [11:0] CSR_SSCRATCHCSW = 12'h148;
  localparam logic [11:0] CSR_SSCRATCHCSWL = 12'h149;
  localparam logic [11:0] CSR_MTVT = 12'h307;
  localparam logic [11:0] CSR_MNXTI = 12'h345;
  localparam logic [11:0] CSR_MINTSTATUS = 12'h346;
  localparam logic [11:0] CSR_MSCRATCHCSW = 12'h348;
  localparam logic [11:0] CSR_MSCRATCHCSWL = 12'h349;
  localparam logic [11:0] CSR_MSTATUS = 12'h300;
  localparam logic [11:0] CSR_MISA = 12'h301;
  localparam logic [11:0] CSR_MEDELEG = 12'h302;
  localparam logic [11:0] CSR_MIDELEG = 12'h303;
  localparam logic [11:0] CSR_MIE = 12'h304;
  localparam logic [11:0] CSR_MTVEC = 12'h305;
  localparam logic [11:0] CSR_MCOUNTEREN = 12'h306;
  localparam logic [11:0] CSR_MSCRATCH = 12'h340;
  localparam logic [11:0] CSR_MEPC = 12'h341;
  localparam logic [11:0] CSR_MCAUSE = 12'h342;
  localparam logic [11:0] CSR_MTVAL = 12'h343;
  localparam logic [11:0] CSR_MIP = 12'h344;
  localparam logic [11:0] CSR_PMPCFG0 = 12'h3a0;
  localparam logic [11:0] CSR_PMPCFG1 = 12'h3a1;
  localparam logic [11:0] CSR_PMPCFG2 = 12'h3a2;
  localparam logic [11:0] CSR_PMPCFG3 = 12'h3a3;
  localparam logic [11:0] CSR_PMPADDR0 = 12'h3b0;
  localparam logic [11:0] CSR_PMPADDR1 = 12'h3b1;
  localparam logic [11:0] CSR_PMPADDR2 = 12'h3b2;
  localparam logic [11:0] CSR_PMPADDR3 = 12'h3b3;
  localparam logic [11:0] CSR_PMPADDR4 = 12'h3b4;
  localparam logic [11:0] CSR_PMPADDR5 = 12'h3b5;
  localparam logic [11:0] CSR_PMPADDR6 = 12'h3b6;
  localparam logic [11:0] CSR_PMPADDR7 = 12'h3b7;
  localparam logic [11:0] CSR_PMPADDR8 = 12'h3b8;
  localparam logic [11:0] CSR_PMPADDR9 = 12'h3b9;
  localparam logic [11:0] CSR_PMPADDR10 = 12'h3ba;
  localparam logic [11:0] CSR_PMPADDR11 = 12'h3bb;
  localparam logic [11:0] CSR_PMPADDR12 = 12'h3bc;
  localparam logic [11:0] CSR_PMPADDR13 = 12'h3bd;
  localparam logic [11:0] CSR_PMPADDR14 = 12'h3be;
  localparam logic [11:0] CSR_PMPADDR15 = 12'h3bf;
  localparam logic [11:0] CSR_TSELECT = 12'h7a0;
  localparam logic [11:0] CSR_TDATA1 = 12'h7a1;
  localparam logic [11:0] CSR_TDATA2 = 12'h7a2;
  localparam logic [11:0] CSR_TDATA3 = 12'h7a3;
  localparam logic [11:0] CSR_DCSR = 12'h7b0;
  localparam logic [11:0] CSR_DPC = 12'h7b1;
  localparam logic [11:0] CSR_DSCRATCH = 12'h7b2;
  localparam logic [11:0] CSR_MCYCLE = 12'hb00;
  localparam logic [11:0] CSR_MINSTRET = 12'hb02;
  localparam logic [11:0] CSR_MHPMCOUNTER3 = 12'hb03;
  localparam logic [11:0] CSR_MHPMCOUNTER4 = 12'hb04;
  localparam logic [11:0] CSR_MHPMCOUNTER5 = 12'hb05;
  localparam logic [11:0] CSR_MHPMCOUNTER6 = 12'hb06;
  localparam logic [11:0] CSR_MHPMCOUNTER7 = 12'hb07;
  localparam logic [11:0] CSR_MHPMCOUNTER8 = 12'hb08;
  localparam logic [11:0] CSR_MHPMCOUNTER9 = 12'hb09;
  localparam logic [11:0] CSR_MHPMCOUNTER10 = 12'hb0a;
  localparam logic [11:0] CSR_MHPMCOUNTER11 = 12'hb0b;
  localparam logic [11:0] CSR_MHPMCOUNTER12 = 12'hb0c;
  localparam logic [11:0] CSR_MHPMCOUNTER13 = 12'hb0d;
  localparam logic [11:0] CSR_MHPMCOUNTER14 = 12'hb0e;
  localparam logic [11:0] CSR_MHPMCOUNTER15 = 12'hb0f;
  localparam logic [11:0] CSR_MHPMCOUNTER16 = 12'hb10;
  localparam logic [11:0] CSR_MHPMCOUNTER17 = 12'hb11;
  localparam logic [11:0] CSR_MHPMCOUNTER18 = 12'hb12;
  localparam logic [11:0] CSR_MHPMCOUNTER19 = 12'hb13;
  localparam logic [11:0] CSR_MHPMCOUNTER20 = 12'hb14;
  localparam logic [11:0] CSR_MHPMCOUNTER21 = 12'hb15;
  localparam logic [11:0] CSR_MHPMCOUNTER22 = 12'hb16;
  localparam logic [11:0] CSR_MHPMCOUNTER23 = 12'hb17;
  localparam logic [11:0] CSR_MHPMCOUNTER24 = 12'hb18;
  localparam logic [11:0] CSR_MHPMCOUNTER25 = 12'hb19;
  localparam logic [11:0] CSR_MHPMCOUNTER26 = 12'hb1a;
  localparam logic [11:0] CSR_MHPMCOUNTER27 = 12'hb1b;
  localparam logic [11:0] CSR_MHPMCOUNTER28 = 12'hb1c;
  localparam logic [11:0] CSR_MHPMCOUNTER29 = 12'hb1d;
  localparam logic [11:0] CSR_MHPMCOUNTER30 = 12'hb1e;
  localparam logic [11:0] CSR_MHPMCOUNTER31 = 12'hb1f;
  localparam logic [11:0] CSR_MHPMEVENT3 = 12'h323;
  localparam logic [11:0] CSR_MHPMEVENT4 = 12'h324;
  localparam logic [11:0] CSR_MHPMEVENT5 = 12'h325;
  localparam logic [11:0] CSR_MHPMEVENT6 = 12'h326;
  localparam logic [11:0] CSR_MHPMEVENT7 = 12'h327;
  localparam logic [11:0] CSR_MHPMEVENT8 = 12'h328;
  localparam logic [11:0] CSR_MHPMEVENT9 = 12'h329;
  localparam logic [11:0] CSR_MHPMEVENT10 = 12'h32a;
  localparam logic [11:0] CSR_MHPMEVENT11 = 12'h32b;
  localparam logic [11:0] CSR_MHPMEVENT12 = 12'h32c;
  localparam logic [11:0] CSR_MHPMEVENT13 = 12'h32d;
  localparam logic [11:0] CSR_MHPMEVENT14 = 12'h32e;
  localparam logic [11:0] CSR_MHPMEVENT15 = 12'h32f;
  localparam logic [11:0] CSR_MHPMEVENT16 = 12'h330;
  localparam logic [11:0] CSR_MHPMEVENT17 = 12'h331;
  localparam logic [11:0] CSR_MHPMEVENT18 = 12'h332;
  localparam logic [11:0] CSR_MHPMEVENT19 = 12'h333;
  localparam logic [11:0] CSR_MHPMEVENT20 = 12'h334;
  localparam logic [11:0] CSR_MHPMEVENT21 = 12'h335;
  localparam logic [11:0] CSR_MHPMEVENT22 = 12'h336;
  localparam logic [11:0] CSR_MHPMEVENT23 = 12'h337;
  localparam logic [11:0] CSR_MHPMEVENT24 = 12'h338;
  localparam logic [11:0] CSR_MHPMEVENT25 = 12'h339;
  localparam logic [11:0] CSR_MHPMEVENT26 = 12'h33a;
  localparam logic [11:0] CSR_MHPMEVENT27 = 12'h33b;
  localparam logic [11:0] CSR_MHPMEVENT28 = 12'h33c;
  localparam logic [11:0] CSR_MHPMEVENT29 = 12'h33d;
  localparam logic [11:0] CSR_MHPMEVENT30 = 12'h33e;
  localparam logic [11:0] CSR_MHPMEVENT31 = 12'h33f;
  localparam logic [11:0] CSR_MVENDORID = 12'hf11;
  localparam logic [11:0] CSR_MARCHID = 12'hf12;
  localparam logic [11:0] CSR_MIMPID = 12'hf13;
  localparam logic [11:0] CSR_MHARTID = 12'hf14;
  localparam logic [11:0] CSR_SSR = 12'h7c0;
  localparam logic [11:0] CSR_FPMODE = 12'h7c1;
  localparam logic [11:0] CSR_CYCLEH = 12'hc80;
  localparam logic [11:0] CSR_TIMEH = 12'hc81;
  localparam logic [11:0] CSR_INSTRETH = 12'hc82;
  localparam logic [11:0] CSR_HPMCOUNTER3H = 12'hc83;
  localparam logic [11:0] CSR_HPMCOUNTER4H = 12'hc84;
  localparam logic [11:0] CSR_HPMCOUNTER5H = 12'hc85;
  localparam logic [11:0] CSR_HPMCOUNTER6H = 12'hc86;
  localparam logic [11:0] CSR_HPMCOUNTER7H = 12'hc87;
  localparam logic [11:0] CSR_HPMCOUNTER8H = 12'hc88;
  localparam logic [11:0] CSR_HPMCOUNTER9H = 12'hc89;
  localparam logic [11:0] CSR_HPMCOUNTER10H = 12'hc8a;
  localparam logic [11:0] CSR_HPMCOUNTER11H = 12'hc8b;
  localparam logic [11:0] CSR_HPMCOUNTER12H = 12'hc8c;
  localparam logic [11:0] CSR_HPMCOUNTER13H = 12'hc8d;
  localparam logic [11:0] CSR_HPMCOUNTER14H = 12'hc8e;
  localparam logic [11:0] CSR_HPMCOUNTER15H = 12'hc8f;
  localparam logic [11:0] CSR_HPMCOUNTER16H = 12'hc90;
  localparam logic [11:0] CSR_HPMCOUNTER17H = 12'hc91;
  localparam logic [11:0] CSR_HPMCOUNTER18H = 12'hc92;
  localparam logic [11:0] CSR_HPMCOUNTER19H = 12'hc93;
  localparam logic [11:0] CSR_HPMCOUNTER20H = 12'hc94;
  localparam logic [11:0] CSR_HPMCOUNTER21H = 12'hc95;
  localparam logic [11:0] CSR_HPMCOUNTER22H = 12'hc96;
  localparam logic [11:0] CSR_HPMCOUNTER23H = 12'hc97;
  localparam logic [11:0] CSR_HPMCOUNTER24H = 12'hc98;
  localparam logic [11:0] CSR_HPMCOUNTER25H = 12'hc99;
  localparam logic [11:0] CSR_HPMCOUNTER26H = 12'hc9a;
  localparam logic [11:0] CSR_HPMCOUNTER27H = 12'hc9b;
  localparam logic [11:0] CSR_HPMCOUNTER28H = 12'hc9c;
  localparam logic [11:0] CSR_HPMCOUNTER29H = 12'hc9d;
  localparam logic [11:0] CSR_HPMCOUNTER30H = 12'hc9e;
  localparam logic [11:0] CSR_HPMCOUNTER31H = 12'hc9f;
  localparam logic [11:0] CSR_MCYCLEH = 12'hb80;
  localparam logic [11:0] CSR_MINSTRETH = 12'hb82;
  localparam logic [11:0] CSR_MHPMCOUNTER3H = 12'hb83;
  localparam logic [11:0] CSR_MHPMCOUNTER4H = 12'hb84;
  localparam logic [11:0] CSR_MHPMCOUNTER5H = 12'hb85;
  localparam logic [11:0] CSR_MHPMCOUNTER6H = 12'hb86;
  localparam logic [11:0] CSR_MHPMCOUNTER7H = 12'hb87;
  localparam logic [11:0] CSR_MHPMCOUNTER8H = 12'hb88;
  localparam logic [11:0] CSR_MHPMCOUNTER9H = 12'hb89;
  localparam logic [11:0] CSR_MHPMCOUNTER10H = 12'hb8a;
  localparam logic [11:0] CSR_MHPMCOUNTER11H = 12'hb8b;
  localparam logic [11:0] CSR_MHPMCOUNTER12H = 12'hb8c;
  localparam logic [11:0] CSR_MHPMCOUNTER13H = 12'hb8d;
  localparam logic [11:0] CSR_MHPMCOUNTER14H = 12'hb8e;
  localparam logic [11:0] CSR_MHPMCOUNTER15H = 12'hb8f;
  localparam logic [11:0] CSR_MHPMCOUNTER16H = 12'hb90;
  localparam logic [11:0] CSR_MHPMCOUNTER17H = 12'hb91;
  localparam logic [11:0] CSR_MHPMCOUNTER18H = 12'hb92;
  localparam logic [11:0] CSR_MHPMCOUNTER19H = 12'hb93;
  localparam logic [11:0] CSR_MHPMCOUNTER20H = 12'hb94;
  localparam logic [11:0] CSR_MHPMCOUNTER21H = 12'hb95;
  localparam logic [11:0] CSR_MHPMCOUNTER22H = 12'hb96;
  localparam logic [11:0] CSR_MHPMCOUNTER23H = 12'hb97;
  localparam logic [11:0] CSR_MHPMCOUNTER24H = 12'hb98;
  localparam logic [11:0] CSR_MHPMCOUNTER25H = 12'hb99;
  localparam logic [11:0] CSR_MHPMCOUNTER26H = 12'hb9a;
  localparam logic [11:0] CSR_MHPMCOUNTER27H = 12'hb9b;
  localparam logic [11:0] CSR_MHPMCOUNTER28H = 12'hb9c;
  localparam logic [11:0] CSR_MHPMCOUNTER29H = 12'hb9d;
  localparam logic [11:0] CSR_MHPMCOUNTER30H = 12'hb9e;
  localparam logic [11:0] CSR_MHPMCOUNTER31H = 12'hb9f;
endpackage
// verilog_lint: waive-stop parameter-name-style
